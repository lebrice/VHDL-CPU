entity fetchStage is
  port (
    clock
  ) ;
end fetchStage;

architecture fetchStage_arch of fetchStage is



begin



end architecture ; -- arch