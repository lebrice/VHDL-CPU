library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity fetchStage is
  port (
    clock : std_logic
  ) ;
end fetchStage;

architecture fetchStage_arch of fetchStage is



begin



end architecture ; -- arch