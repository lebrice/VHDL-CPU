entity memoryStage is
  port (
    clock
  ) ;
end memoryStage ;

architecture memoryStage_arch of memoryStage is



begin



end architecture ; -- arch