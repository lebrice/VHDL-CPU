entity decodeStage is
  port (
    clock
  ) ;
end decodeStage ;

architecture decodeStage_arch of decodeStage is



begin



end architecture ; -- arch