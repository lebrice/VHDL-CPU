library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity memoryStage is
  port (
    clock : in std_logic;
  ) ;
end memoryStage ;

architecture memoryStage_arch of memoryStage is



begin



end architecture ; -- arch