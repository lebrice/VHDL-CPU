library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity decodeStage is
  port (
    clock : std_logic
  ) ;
end decodeStage ;

architecture decodeStage_arch of decodeStage is



begin



end architecture ; -- arch