library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity writebackStage is
  port (
    clock : std_logic
  ) ;
end writebackStage ;

architecture writebackStage_arch of writebackStage is



begin



end architecture ; -- arch