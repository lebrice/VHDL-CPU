entity executeStage is
  port (
    clock
  ) ;
end executeStage ;

architecture executeStage_arch of executeStage is



begin



end architecture ; -- arch