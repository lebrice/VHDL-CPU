library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity executeStage is
  port (
    clock : std_logic
  ) ;
end executeStage ;

architecture executeStage_arch of executeStage is



begin



end architecture ; -- arch