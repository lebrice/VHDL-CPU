library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_textio.all;
    use ieee.numeric_std.all;


    package fifo is

    end fifo;

    package body fifo is

    end fifo;