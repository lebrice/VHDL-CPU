entity ALU is
  port (
    clock
  ) ;
end ALU ;

architecture ALU_arch of ALU is



begin



end architecture ; -- arch