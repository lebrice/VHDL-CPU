library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity processor is
  port (
    clock : std_logic
  ) ;
end processor;

architecture pipeline_processor_arch of processor is



begin



end architecture ; -- arch