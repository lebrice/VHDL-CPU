entity processor is
  port (
    clock
  ) ;
end processor;

architecture pipeline_processor_arch of processor is



begin



end architecture ; -- arch